module cpu (
    input  wire        clk,
    input  wire        rst,
    input  logic [31:0] instruction_in, // direct instruction feed for testing

    output logic [31:0] readd // observation signal for testing
);


/*
my thoughts but wires for lw instruction

GETTING DATA MEMORY
read_data from data                     -> write_data for registers
    alu_add(rs1+sign extended immediate)    -> read_data_adress (data_memory in port)
    read_data                               -> data_memory (adress in port([31:0]) write_data out port([31:0]))

WRITING TO REGISTERS
destination_register(control out port)  -> register_adress (regfile in port)
reg_write (control out port)            -> enabled ()

decoder -> control


*/


// WIRES BETWEEN COMPONENTS NOT FROM INSTRUCTIONS
logic [31:0] regData; // unused placeholder for future instructions
logic [31:0] dData; // out from data memory, in to reg file
logic [3:0]  alu_ctrl; // control word into ALU
logic [31:0] data_address; // data address to be read (wire between the ALU out and the data memory)
logic        reg_write; // 1 bit wire from control to registers
logic [3:0]  inst_type;
logic [2:0]  imm_type; // used only by the sign extender
logic [31:0] regData1;
logic [31:0] regData2;
logic        memRead;
logic        memWrite;
logic        alu_zero;
logic        alu_last_bit;

// WIRES DIRECTLY FROM INSTRUCTION
logic [31:0] instruction;
logic [4:0] rs1;
logic [4:0] rs2;
logic [31:0] immediate;
logic [6:0] opcode;
logic [2:0] func3;
logic [6:0] func7;
logic [4:0] rd;
logic [4:0] reg_destination;
// NEW BUS DLC COMING SOON*tm*




// initiats the program counter as a single register, then counts up (ignore this for the time being, I cant count a program if I cant add generally, this is a placeholder anyway)
                    // reg [31:0] pc;
                    // logic [31:0] next_pc;

                    // always_comb begin : pcSelect
                    //     next_pc = pc + 4; // forward 4 bits
                    // end

                    // // zeros the program counter when done 
                    // always @(posedge clk) begin
                    //     if (rst = 0)
                    //         pc = 32'b0; 
                    // end







// memory #(
//     .mem_init("") // file path to ADD ONCE I HAVE A FILE  ignore this for now :)
// ) instruction_memory (
//     // Memory inputs
//     .clk(clk), // Connects clk of each module to higher level speficied port (weird module hierarchy thing)
//     .address(pc),
//     .write_data(32'b0), // when nothing to connect to, im defining them as wires of the correct width
//     .write_enable(1'b0),
//     .rst_n(1'b1),

//     // Memory outputs
//     .read_data(instruction)
// );

// Register File
registerFile register_file_inst (
    .clk(clk),
    .rst(rst),
    .rs1(rs1),
    .rs2(rs2),
    .rd(reg_destination),
    .wd(dData),
    .enableWrite(reg_write),
    .rd1(regData1),
    .rd2(regData2)
);

// Data Memory
dataMemory data_memory_inst (
    .clk(clk),
    .address(data_address),
    .write_data(regData2),
    .write_enable(memWrite),
    .rst_data(rst),
    .read_data(dData)
);

<<<<<<< HEAD
<<<<<<< HEAD
// ALU for data memory adress calculation
alu (
    .clk(clk)
    .rst(rst)
    .cntrl(alu_op) // from control module, control must be modified further to support different functions per inst type
    .d1(regData1)
    .d2(immediate)                      // MAKE THIS THE SIGN EXTENDED IMMEDIATE 

    .alu_output(data_adress) // to data memory
    .zero                               // useless ports, I already know what zero is im sure the machine can do the same
    .last_bit
)
=======
=======
>>>>>>> b9e8ade2a854973ddec0436419768f4e07dc0613
// ALU for data memory address calculation
alu alu_inst (
    .clk(clk),
    .rst(rst),
    .cntrl(alu_ctrl),
    .d1(regData1),
    .d2(immediate),
    .alu_output(data_address),
    .zero(alu_zero),
    .last_bit(alu_last_bit)
);
<<<<<<< HEAD
>>>>>>> b9e8ade2a854973ddec0436419768f4e07dc0613
=======
>>>>>>> b9e8ade2a854973ddec0436419768f4e07dc0613

// Control unit
control control_inst (
    .op(opcode),
    .func3(func3),
    .func7(func7),
    .alu_zero(alu_zero),
    .alu_last_bit(alu_last_bit),
    .alu_control(),
    .imm_source(),
    .mem_read(memRead),
    .mem_write(memWrite),
    .reg_write(reg_write),
    .alu_source(),
    .pc_source(),
    .alu_op(alu_ctrl)
);

// Sign extender
signExtender sign_extender_inst (
    .clk(clk),
    .rst(rst),
    .inst(instruction),
    .imm_type(imm_type),
    .ext_imm(immediate)
);

// Decoder
decoder decoder_inst (
    .clk(clk),
    .rst(rst),
    .instruction(instruction),
    .inst_type(inst_type),
    .rd(reg_destination),
    .rs1(rs1),
    .rs2(rs2),
    .func3(func3),
    .func7(func7),
    .imm_type(imm_type),
    .opcode(opcode),
    .immediate()
);

// direct instruction drive for this testbench-style hookup
assign instruction = instruction_in;

// expose loaded data for visibility
assign readd = dData;

endmodule